// This is a single line comment
// module main
/*
	This is a multi line comment
	/* It can even be nested. */
*/

fn main() {
	println('Hello World')	
}
